
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity RAM32_b is
end RAM32_b;

architecture Behavioral of RAM32_b is

begin


end Behavioral;

