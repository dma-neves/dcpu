

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ROM is
Port(
	adr : in STD_LOGIC_VECTOR(15 downto 0);
	En : in STD_LOGIC;
	DO : out STD_LOGIC_VECTOR(15 downto 0)
);
end ROM;

architecture Behavioral of ROM is

begin

process(adr, En)
begin

	if En = '0' then
		DO <= "0000000000000000";
	else
		
		case adr is
            when "0000000000000000" => DO <= "0000000000010011";
            when "0000000000000001" => DO <= "0000000010000111";
            when "0000000000000010" => DO <= "0000000000000100";
            when "0000000000000011" => DO <= "0000000000000111";
            when "0000000000000100" => DO <= "0000000000001110";
            when "0000000000000101" => DO <= "0000000000000111";
            when "0000000000000110" => DO <= "0000000000001101";
            when "0000000000000111" => DO <= "0000000000000111";
            when "0000000000001000" => DO <= "0000000000001011";
            when "0000000000001001" => DO <= "0000000000000001";
            when "0000000000001010" => DO <= "0000000000000100";
            when "0000000000001011" => DO <= "0000000000000111";
            when "0000000000001100" => DO <= "0000000000001110";
            when "0000000000001101" => DO <= "0000000000000111";
            when "0000000000001110" => DO <= "0000000000001101";
            when "0000000000001111" => DO <= "0000000000000111";
            when "0000000000010000" => DO <= "0000000000001011";
            when "0000000000010001" => DO <= "0000000000000010";
            when "0000000000010010" => DO <= "0000000000001001";
            when "0000000000010011" => DO <= "0000000000111110";
            when "0000000000010100" => DO <= "0000000000001010";
            when "0000000000010101" => DO <= "0000000000000000";
            when "0000000000010110" => DO <= "0000000000001011";
            when "0000000000010111" => DO <= "0000000000000011";
            when "0000000000011000" => DO <= "0000000000001001";
            when "0000000000011001" => DO <= "0000000000111110";
            when "0000000000011010" => DO <= "0000000000001010";
            when "0000000000011011" => DO <= "0000000000000000";
            when "0000000000011100" => DO <= "0000000000001011";
            when "0000000000011101" => DO <= "0000000000000100";
            when "0000000000011110" => DO <= "0000000000000001";
            when "0000000000011111" => DO <= "0000010000000010";
            when "0000000000100000" => DO <= "0000000000010101";
            when "0000000000100001" => DO <= "0000000000110011";
            when "0000000000100010" => DO <= "0000000000010100";
            when "0000000000100011" => DO <= "0000000000110011";
            when "0000000000100100" => DO <= "0000000000000000";
            when "0000000000100101" => DO <= "0000010000000001";
            when "0000000000100110" => DO <= "0000000000001111";
            when "0000000000100111" => DO <= "0000000000000000";
            when "0000000000101000" => DO <= "0000000000001011";
            when "0000000000101001" => DO <= "0000000000000101";
            when "0000000000101010" => DO <= "0000000000000000";
            when "0000000000101011" => DO <= "0000010100000011";
            when "0000000000101100" => DO <= "0000000000001110";
            when "0000000000101101" => DO <= "0000000000000011";
            when "0000000000101110" => DO <= "0000000000000011";
            when "0000000000101111" => DO <= "0000000000000100";
            when "0000000000110000" => DO <= "0000000000001110";
            when "0000000000110001" => DO <= "0000000000000100";
            when "0000000000110010" => DO <= "0000000000010011";
            when "0000000000110011" => DO <= "0000000000011101";
            when "0000000000110100" => DO <= "0000000000001101";
            when "0000000000110101" => DO <= "0000000000000111";
            when "0000000000110110" => DO <= "0000000000001010";
            when "0000000000110111" => DO <= "0000000000000000";
            when "0000000000111000" => DO <= "0000000000000011";
            when "0000000000111001" => DO <= "0000000000000111";
            when "0000000000111010" => DO <= "0000000000001110";
            when "0000000000111011" => DO <= "0000000000000111";
            when "0000000000111100" => DO <= "0000000000001101";
            when "0000000000111101" => DO <= "0000000000000111";
            when "0000000000111110" => DO <= "0000000000001100";
            when "0000000000111111" => DO <= "0000000000000011";
            when "0000000001000000" => DO <= "0000000000000011";
            when "0000000001000001" => DO <= "0000000000000111";
            when "0000000001000010" => DO <= "0000000000001110";
            when "0000000001000011" => DO <= "0000000000000111";
            when "0000000001000100" => DO <= "0000000000000010";
            when "0000000001000101" => DO <= "0000000000000001";
            when "0000000001000110" => DO <= "0000000000001111";
            when "0000000001000111" => DO <= "0000000000000000";
            when "0000000001001000" => DO <= "0000000000001011";
            when "0000000001001001" => DO <= "0000000000000101";
            when "0000000001001010" => DO <= "0000000000000001";
            when "0000000001001011" => DO <= "0000001000000101";
            when "0000000001001100" => DO <= "0000000000001110";
            when "0000000001001101" => DO <= "0000000000000101";
            when "0000000001001110" => DO <= "0000000000000010";
            when "0000000001001111" => DO <= "0000000000000001";
            when "0000000001010000" => DO <= "0000000000001111";
            when "0000000001010001" => DO <= "0000000000000000";
            when "0000000001010010" => DO <= "0000000000001100";
            when "0000000001010011" => DO <= "0000000000000101";
            when "0000000001010100" => DO <= "0000000000000010";
            when "0000000001010101" => DO <= "0000000000000001";
            when "0000000001010110" => DO <= "0000000000001111";
            when "0000000001010111" => DO <= "0000000000000000";
            when "0000000001011000" => DO <= "0000000000001011";
            when "0000000001011001" => DO <= "0000000000000101";
            when "0000000001011010" => DO <= "0000000000000100";
            when "0000000001011011" => DO <= "0000000000000101";
            when "0000000001011100" => DO <= "0000000000010101";
            when "0000000001011101" => DO <= "0000000001101111";
            when "0000000001011110" => DO <= "0000000000000010";
            when "0000000001011111" => DO <= "0000000000000010";
            when "0000000001100000" => DO <= "0000000000001111";
            when "0000000001100001" => DO <= "0000000000000000";
            when "0000000001100010" => DO <= "0000000000001011";
            when "0000000001100011" => DO <= "0000000000000101";
            when "0000000001100100" => DO <= "0000000000000011";
            when "0000000001100101" => DO <= "0000000000000101";
            when "0000000001100110" => DO <= "0000000000001110";
            when "0000000001100111" => DO <= "0000000000000101";
            when "0000000001101000" => DO <= "0000000000000010";
            when "0000000001101001" => DO <= "0000000000000010";
            when "0000000001101010" => DO <= "0000000000001111";
            when "0000000001101011" => DO <= "0000000000000000";
            when "0000000001101100" => DO <= "0000000000001100";
            when "0000000001101101" => DO <= "0000000000000101";
            when "0000000001101110" => DO <= "0000000000010011";
            when "0000000001101111" => DO <= "0000000001000011";
            when "0000000001110000" => DO <= "0000000000000100";
            when "0000000001110001" => DO <= "0000000000000111";
            when "0000000001110010" => DO <= "0000000000001110";
            when "0000000001110011" => DO <= "0000000000000111";
            when "0000000001110100" => DO <= "0000000000000100";
            when "0000000001110101" => DO <= "0000000000000111";
            when "0000000001110110" => DO <= "0000000000001110";
            when "0000000001110111" => DO <= "0000000000000111";
            when "0000000001111000" => DO <= "0000000000001101";
            when "0000000001111001" => DO <= "0000000000000111";
            when "0000000001111010" => DO <= "0000000000001011";
            when "0000000001111011" => DO <= "0000000000000000";
            when "0000000001111100" => DO <= "0000000000000100";
            when "0000000001111101" => DO <= "0000000000000111";
            when "0000000001111110" => DO <= "0000000000001110";
            when "0000000001111111" => DO <= "0000000000000111";
            when "0000000010000000" => DO <= "0000000000001101";
            when "0000000010000001" => DO <= "0000000000000111";
            when "0000000010000010" => DO <= "0000000000001011";
            when "0000000010000011" => DO <= "0000000000000001";
            when "0000000010000100" => DO <= "0000000000001101";
            when "0000000010000101" => DO <= "0000000000000001";
            when "0000000010000110" => DO <= "0000000000010010";
            when "0000000010000111" => DO <= "0000000000000000";
            when "0000000010001000" => DO <= "0000000000001101";
            when "0000000010001001" => DO <= "0000000000000111";
            when "0000000010001010" => DO <= "0000000000001010";
            when "0000000010001011" => DO <= "0000000000000011";
            when "0000000010001100" => DO <= "0000000000000011";
            when "0000000010001101" => DO <= "0000000000000111";
            when "0000000010001110" => DO <= "0000000000001110";
            when "0000000010001111" => DO <= "0000000000000111";
            when "0000000010010000" => DO <= "0000000000001101";
            when "0000000010010001" => DO <= "0000000000000111";
            when "0000000010010010" => DO <= "0000000000001010";
            when "0000000010010011" => DO <= "0000000000000101";
            when "0000000010010100" => DO <= "0000000000000011";
            when "0000000010010101" => DO <= "0000000000000111";
            when "0000000010010110" => DO <= "0000000000001110";
            when "0000000010010111" => DO <= "0000000000000111";
            when "0000000010011000" => DO <= "0000000000001101";
            when "0000000010011001" => DO <= "0000000000000111";
            when "0000000010011010" => DO <= "0000000000001010";
            when "0000000010011011" => DO <= "0000000000000010";
            when "0000000010011100" => DO <= "0000000000000011";
            when "0000000010011101" => DO <= "0000000000000111";
            when "0000000010011110" => DO <= "0000000000001110";
            when "0000000010011111" => DO <= "0000000000000111";
            when "0000000010100000" => DO <= "0000000000001101";
            when "0000000010100001" => DO <= "0000000000000111";
            when "0000000010100010" => DO <= "0000000000001010";
            when "0000000010100011" => DO <= "0000000000001001";
            when "0000000010100100" => DO <= "0000000000000011";
            when "0000000010100101" => DO <= "0000000000000111";
            when "0000000010100110" => DO <= "0000000000001110";
            when "0000000010100111" => DO <= "0000000000000111";
            when "0000000010101000" => DO <= "0000000000001101";
            when "0000000010101001" => DO <= "0000000000000111";
            when "0000000010101010" => DO <= "0000000000001010";
            when "0000000010101011" => DO <= "0000000011001001";
            when "0000000010101100" => DO <= "0000000000000011";
            when "0000000010101101" => DO <= "0000000000000111";
            when "0000000010101110" => DO <= "0000000000001110";
            when "0000000010101111" => DO <= "0000000000000111";
            when "0000000010110000" => DO <= "0000000000000010";
            when "0000000010110001" => DO <= "0000000000000101";
            when "0000000010110010" => DO <= "0000000000001111";
            when "0000000010110011" => DO <= "0000000000000000";
            when "0000000010110100" => DO <= "0000000000001011";
            when "0000000010110101" => DO <= "0000000000000000";
            when "0000000010110110" => DO <= "0000000000001101";
            when "0000000010110111" => DO <= "0000000000000111";
            when "0000000010111000" => DO <= "0000000000001100";
            when "0000000010111001" => DO <= "0000000000000000";
            when "0000000010111010" => DO <= "0000000000000011";
            when "0000000010111011" => DO <= "0000000000000111";
            when "0000000010111100" => DO <= "0000000000001110";
            when "0000000010111101" => DO <= "0000000000000111";
            when "0000000010111110" => DO <= "0000000000000010";
            when "0000000010111111" => DO <= "0000000000000101";
            when "0000000011000000" => DO <= "0000000000001101";
            when "0000000011000001" => DO <= "0000000000000111";
            when "0000000011000010" => DO <= "0000000000010000";
            when "0000000011000011" => DO <= "0000000000000000";
            when "0000000011000100" => DO <= "0000000000000011";
            when "0000000011000101" => DO <= "0000000000000111";
            when "0000000011000110" => DO <= "0000000000001110";
            when "0000000011000111" => DO <= "0000000000000111";
            when "0000000011001000" => DO <= "0000000000010011";
            when "0000000011001001" => DO <= "0000000000000001";
            when "0000000011001010" => DO <= "0000000000010111";
            when "0000000011001011" => DO <= "0000000000000000";

            when others => DO <= "0000000000000000";
		end case;
		
	end if;

end process;

end Behavioral;
